`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Student: Tawseef Patel 101145333 & Saad Babur 101123210
// 
// Create Date: 10/14/2022
// Design Name: lab1_2_1.v 
// Module Name: lab1_2_1
// Project Name: Lab 1_2
//////////////////////////////////////////////////////////////////////////////////


module lab1_2_1(
    input [7:0]x_in,
    output [7:0]y_out
    );
    
    assign y_out = x_in;
    
endmodule
