`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Student: Tawseef Patel 101145333 & Saad Babur 101123210
// 
// Create Date: 10/14/2022 03:41:20 PM
// Design Name: 2x1 MUX - GATE LEVEL 
// Module Name: lab1_1_1
// Project Name: Lab 1
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module lab1_2_1(
    input [7:0]x_in,
    output [7:0]y_out
    );
    
    assign y_out = x_in;
    
endmodule
